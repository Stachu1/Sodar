library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sodar_ip_v1_0 is
	generic (
        DUTY_DEFAULT    : std_logic_vector(31 downto 0) := x"000000C8";  -- Example: decimal 200
        PERIOD_DEFAULT  : std_logic_vector(31 downto 0) := x"00000190";  -- Example: decimal 400
        PHASE_DEFAULT   : std_logic_vector(31 downto 0) := x"00000003";


		-- Parameters of Axi Slave Bus Interface S00_AXI
		C_S00_AXI_DATA_WIDTH	: integer	:= 32;
		C_S00_AXI_ADDR_WIDTH	: integer	:= 4
	);
	port (
		-- Users to add ports here

		-- User ports ends
		-- Do not modify the ports beyond this line
        duty_cycle : out std_logic_vector(C_S00_AXI_DATA_WIDTH-1 downto 0);
        period     : out std_logic_vector(C_S00_AXI_DATA_WIDTH-1 downto 0);
        phase      : out std_logic_vector(C_S00_AXI_DATA_WIDTH-1 downto 0);

		-- Ports of Axi Slave Bus Interface S00_AXI
		s00_axi_aclk	: in std_logic;
		s00_axi_aresetn	: in std_logic;
		s00_axi_awaddr	: in std_logic_vector(C_S00_AXI_ADDR_WIDTH-1 downto 0);
		s00_axi_awprot	: in std_logic_vector(2 downto 0);
		s00_axi_awvalid	: in std_logic;
		s00_axi_awready	: out std_logic;
		s00_axi_wdata	: in std_logic_vector(C_S00_AXI_DATA_WIDTH-1 downto 0);
		s00_axi_wstrb	: in std_logic_vector((C_S00_AXI_DATA_WIDTH/8)-1 downto 0);
		s00_axi_wvalid	: in std_logic;
		s00_axi_wready	: out std_logic;
		s00_axi_bresp	: out std_logic_vector(1 downto 0);
		s00_axi_bvalid	: out std_logic;
		s00_axi_bready	: in std_logic;
		s00_axi_araddr	: in std_logic_vector(C_S00_AXI_ADDR_WIDTH-1 downto 0);
		s00_axi_arprot	: in std_logic_vector(2 downto 0);
		s00_axi_arvalid	: in std_logic;
		s00_axi_arready	: out std_logic;
		s00_axi_rdata	: out std_logic_vector(C_S00_AXI_DATA_WIDTH-1 downto 0);
		s00_axi_rresp	: out std_logic_vector(1 downto 0);
		s00_axi_rvalid	: out std_logic;
		s00_axi_rready	: in std_logic
	);
end sodar_ip_v1_0;

architecture arch_imp of sodar_ip_v1_0 is

	-- component declaration
	component sodar_ip_v1_0_S00_AXI is
		generic (
		C_S_AXI_DATA_WIDTH	: integer	:= 32;
		C_S_AXI_ADDR_WIDTH	: integer	:= 4
		);
		port (
		S_AXI_ACLK	: in std_logic;
		S_AXI_ARESETN	: in std_logic;
		S_AXI_AWADDR	: in std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
		S_AXI_AWPROT	: in std_logic_vector(2 downto 0);
		S_AXI_AWVALID	: in std_logic;
		S_AXI_AWREADY	: out std_logic;
		S_AXI_WDATA	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
		S_AXI_WSTRB	: in std_logic_vector((C_S_AXI_DATA_WIDTH/8)-1 downto 0);
		S_AXI_WVALID	: in std_logic;
		S_AXI_WREADY	: out std_logic;
		S_AXI_BRESP	: out std_logic_vector(1 downto 0);
		S_AXI_BVALID	: out std_logic;
		S_AXI_BREADY	: in std_logic;
		S_AXI_ARADDR	: in std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
		S_AXI_ARPROT	: in std_logic_vector(2 downto 0);
		S_AXI_ARVALID	: in std_logic;
		S_AXI_ARREADY	: out std_logic;
		S_AXI_RDATA	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
		S_AXI_RRESP	: out std_logic_vector(1 downto 0);
		S_AXI_RVALID	: out std_logic;
		S_AXI_RREADY	: in std_logic
		);
	end component sodar_ip_v1_0_S00_AXI;
    
    signal reg_duty   : std_logic_vector(C_S00_AXI_DATA_WIDTH-1 downto 0);
    signal reg_period : std_logic_vector(C_S00_AXI_DATA_WIDTH-1 downto 0);
    signal reg_phase  : std_logic_vector(C_S00_AXI_DATA_WIDTH-1 downto 0);
    
begin

-- Instantiation of Axi Bus Interface S00_AXI
sodar_ip_v1_0_S00_AXI_inst : sodar_ip_v1_0_S00_AXI
	generic map (
		C_S_AXI_DATA_WIDTH	=> C_S00_AXI_DATA_WIDTH,
		C_S_AXI_ADDR_WIDTH	=> C_S00_AXI_ADDR_WIDTH
	)
	port map (
		S_AXI_ACLK	=> s00_axi_aclk,
		S_AXI_ARESETN	=> s00_axi_aresetn,
		S_AXI_AWADDR	=> s00_axi_awaddr,
		S_AXI_AWPROT	=> s00_axi_awprot,
		S_AXI_AWVALID	=> s00_axi_awvalid,
		S_AXI_AWREADY	=> s00_axi_awready,
		S_AXI_WDATA	=> s00_axi_wdata,
		S_AXI_WSTRB	=> s00_axi_wstrb,
		S_AXI_WVALID	=> s00_axi_wvalid,
		S_AXI_WREADY	=> s00_axi_wready,
		S_AXI_BRESP	=> s00_axi_bresp,
		S_AXI_BVALID	=> s00_axi_bvalid,
		S_AXI_BREADY	=> s00_axi_bready,
		S_AXI_ARADDR	=> s00_axi_araddr,
		S_AXI_ARPROT	=> s00_axi_arprot,
		S_AXI_ARVALID	=> s00_axi_arvalid,
		S_AXI_ARREADY	=> s00_axi_arready,
		S_AXI_RDATA	=> s00_axi_rdata,
		S_AXI_RRESP	=> s00_axi_rresp,
		S_AXI_RVALID	=> s00_axi_rvalid,
		S_AXI_RREADY	=> s00_axi_rready
	);

	-- Add user logic here
     process(s00_axi_aclk)
        begin
            if rising_edge(s00_axi_aclk) then
                if s00_axi_aresetn = '0' then
                    reg_period <= PERIOD_DEFAULT;
                    reg_duty   <= DUTY_DEFAULT;
                    reg_phase  <= PHASE_DEFAULT;
                else
                    if (s00_axi_awvalid = '1' and s00_axi_wvalid = '1') then
                        case s00_axi_awaddr(3 downto 2) is
                            when "00" =>
                                reg_period <= s00_axi_wdata;
                            when "01" =>
                                reg_duty <= s00_axi_wdata;
                            when "10" =>
                                reg_phase <= s00_axi_wdata;  -- relative phase increment
                            when others =>
                                null;
                        end case;
                    end if;
                end if;
            end if;
        end process;
    
        -- Drive the output ports to be consumed by your PWM generator or top-level PWM module.
        duty_cycle <= reg_duty;
        period     <= reg_period;
        phase      <= reg_phase;
	-- User logic ends

end arch_imp;
